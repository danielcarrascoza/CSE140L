Robertson 

    11111001		   -7 * -6 = 42
   	    1010

    00000000
    1111001 
    000000
-   11001


   00000000						 0000	    1010
   1111001						 11001		 101
   000000						 111001		  10
   00110						 0101010	(-)1
_______1__						 00101010
   00101010  = 42




  101010
																		 -00000000
																		  11111111
	pos * pos multiplier													 +	 1
																		  00000000

        1001		   +9 * 10 = 90
   	    1010													      000000000000
																	  111111111111
																				 1
        1001														 1000000000000
		1010
______________
						0000 1010
		0000			0000 0101
	   1001				1010 0010
	  0000				0101 0001
	 1001
	 1011010


    00001001										e = a+b+c+d
	                 f=0+a
	                 f=f+b
					 f=f+c
					 f=f+d



